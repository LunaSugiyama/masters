// instruction_memory.v
// 命令メモリ (ROMとして実装)

module instruction_memory (
    input wire [31:0] addr,
    output wire [31:0] instruction_out
);

    // 1024ワード (4KB) のメモリを想定
    reg [31:0] mem [0:1023];

    initial begin
        // テスト用の命令
        // I命令:add
        // 例: addi x1, x0, 1  (0x00100093)
        //     addi x2, x0, 2  (0x00200113)
        //     add x3, x1, x2  (0x002081B3)
        //     sub x4, x3, x1  (0x40118233)
        // アドレスはワードアドレス（バイトアドレス/4）で指定
        // mem[0] = 32'h00100093; // addi x1, x0, 1
        // mem[1] = 32'h00200113; // addi x2, x0, 2
        // mem[2] = 32'h002081B3; // add x3, x1, x2 (x3 = x1 + x2 = 1 + 2 = 3)
        // mem[3] = 32'h40118233; // sub x4, x3, x1 (x4 = x3 - x1 = 3 - 1 = 2)

        // テスト用の命令 [funct7][rs2][rs1][funct3][rd][opcode]
       // I-type
        mem[0]  = 32'b000000000001_00000_000_00001_0010011; // addi x1, x0, 1     → x1 = 1
        mem[1]  = 32'b000000000010_00000_000_00010_0010011; // addi x2, x0, 2     → x2 = 2

        // R-type
        mem[2]  = 32'b0000000_00010_00001_000_00011_0110011; // add x3, x1, x2    → x3 = x1 + x2 = 3
        mem[3]  = 32'b0100000_00001_00011_000_00100_0110011; // sub x4, x3, x1    → x4 = x3 - x1 = 2
        mem[4]  = 32'b0000000_00010_00011_100_00101_0110011; // xor x5, x3, x2    → x5 = x3 ^ x2 = 1
        mem[5]  = 32'b0000000_00010_00011_110_00110_0110011; // or  x6, x3, x2    → x6 = x3 | x2 = 3
        mem[6]  = 32'b0000000_00010_00011_111_00111_0110011; // and x7, x3, x2    → x7 = x3 & x2 = 2
        mem[7]  = 32'b0000000_00010_00011_001_01000_0110011; // sll x8, x3, x2    → x8 = x3 << x2 = 12
        mem[8]  = 32'b0000000_00010_00011_101_01001_0110011; // srl x9, x3, x2    → x9 = x3 >> x2 = 0

        // I-type (load, shift)
        // mem[8]  = 32'b000000000000_00010_111_00101_0000011;  // lw   x5, 0(x8)      → x5 = MEM[x8+0]
        // mem[4] = 32'b000000000010_00001_001_01000_0010011;  // slli x8, x1, 2    → x8 = x1 << 2 = 4
        // mem[5] = 32'b010000000010_00001_101_01001_0010011;  // srai x9, x1, 2    → x9 = x1 >>> 2 = 0

        // // S-type
        // mem[5] = 32'b0000000_00101_00010_010_00100_0100011; // sw   x5, 4(x2)      → MEM[x2+0] = x5
        // mem[6] = 32'b000000000100_00010_010_00110_0000011;  // lw   x6, 4(x2)      → x6 = MEM[x2+4]

        // B-type
        // mem[5] = 32'b0000000_00011_00010_000_01000_1100011; // beq x2, x3, +8    → branch not taken
        // mem[6] = 32'b0000000_00011_00010_001_01000_1100011; // bne x2, x3, +8    → branch taken

        // // U-type
        // mem[7] = 32'b00000000000000000001_00101_0110111;   // lui x5, 0x0       → x5 = 0x00000000
        // mem[8] = 32'b00010010001101000101_00001_0110111;   // lui x1, 0x12345  → x13 = 0x12345000

        // // J-type
        // mem[5] = 32'h002000ef;  // jal x1, 4
    end

    assign instruction_out = mem[addr[31:2]]; // バイトアドレスからワードアドレスに変換

endmodule